pBAV       0| �� 1 " k@  �����n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ���������n@   ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    ��������  �n    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ��Ѐ��   � � � � @% %%      ������   � � � � (< <<      ��Ѐ��  	 � � � � 2> >>      ��Ѐ��  
 � � � � FS SS      ��Ѐ��   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � 6O      ��Ѐ�_  � � � � <JN      ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,7  :      �����_  � � � � @< ;A      �����_  � � � � TC B      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  $      �����_  � � � �  r$
       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 6<  @    �����_  � � � � @C AF    �����_  � � � � JH G    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <H  L      �����_  � � � � DO M      ��Ѐ�_  � � � � dnH L      �����_  � � � � dOM      ��Й�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,C        �����_  � � � � dTC       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <<  @    �����_  � � � � DC A    �����_  � � � � dd< @    �����_  � � � � dCA    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        �����_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � C  G      �����_
  � � � � O H      �����_
  � � � � d|C G      �����_
  � � � � d|OH      �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � 7C      �����_  � � � � ddC     ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,T D      �����_  � � � � hT
D    �����_  � � � � T< C      ��У�_  � � � � < C    ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H G    �����_   � � � � @C  F    �����_ ! � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � $        �����_ " � � � � |$       �����_ " � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b���| �J� f T \�Tf�*�X��� ��� 4p � .�                                                                                                                                                                                                                                                                                                                                                                                                                                                          