pBAV        �  ��   @  ����  @   ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������
 @          �����   � � � � 
 @       �����   � � � � 
 @       �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   `D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        