pBAV       �d ��   r@  ����	<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������<@   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������F, $$      ����,�   � � � � h-      �� �	@   � � � � R* **      ����
K   � � � � Z\) ))      ������   � � � � Z$( ((      ������   � � � � ZA1 33      �����_   � � � � Z<2 44      ������   � � � � ZJ3 55      ������   � � � � Z,4 66      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �  @)     �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @F:     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��z�j� 	 � � � �               �����   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O
N      ����+�  � � � � @Dx M      ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ����� 	 � � � � @H      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O
N      ����+�  � � � � @Dx M      ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � H       ������ 
 � � � � @H       ����l� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n@Y       ��ˋl�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 2@Yu       ��ˋl�	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @>       ���O
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @>       ���O  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   vFH�H2����F��\�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              