pBAV       �b ��
   o?  ����
�@?   ���������@?   ���������@?   ���������@?   ���������@?   ���������@?   ���������@?   ���������@?   ���������@?   ���������@?   ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    ��������  �@    �������� b@0 22      ������   � � � �  }@2 33      ������   � � � � uJ- //      ������   � � � � z<2 00      ������   � � � � {,= 11      ������   � � � � ZT) )*      ������   � � � � eT+ ++      ������   � � � �  cT,(--      ������   � � � � g(& &&      ������   � � � � gX" $$      ������   � � � �               ������    � � � �               ������    � � � �               ������    � � � �               ��        � � � �               ��        � � � �               ��        � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I       ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dx     ������ 
 � � � �               ������   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @;0       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T       �����N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @5        ��ڀO  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @D       ��ɀ(�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @P       ����P  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � M@Do     ������	 
 � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �   v����F�	:*\x�H��6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              