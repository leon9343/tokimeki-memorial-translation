pBAV       �  ��   @  �����>?   ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  @$j      �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            