pBAV        � ��   @  �����z@   ���������z@   ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  �z    ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   @:         �����   � � � �   @< $$      �����   � � � �   @@ ((      �����   � � � �   @HF,,      �����   � � � �   @H 00      �����   � � � �   @PF44      �����   � � � �   @P 88      �����   � � � �   @T <<      �����   � � � �   @X @@      �����  	 � � � �   @\ DD      �����  
 � � � �   @` HH      �����   � � � �   @d LL      �����   � � � �   @h PP      �����   � � � �   @0       �����  � � � �   @4       �����  � � � �   @8         �����  � � � �   @< $$      �����  � � � �   @@ ((      �����  � � � �   @D ,,      �����  � � � �   @H 00      �����  � � � �   @L 44      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   � 0pJ2�� h�HD\��6L��8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  