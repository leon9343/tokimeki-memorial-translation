pBAV         ��   @  ����Ʋ@   ��������Ʋ@   ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  Ʋ    ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   r@ ((      �����   � � � �   @; ,,      �����   � � � �   @H 00      �����   � � � �   @L 44      �����   � � � �   @R 88      �����   � � � �   @Y <<      �����  	 � � � �   @^m@@      �����  
 � � � �   @\ DD      �����   � � � �   h HH      �����   � � � �   @m LL      �����  	 � � � �   A ((      �����   � � � �   |g HH      �����   � � � �   @< $$      �����   � � � �   @0       �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   J�d~�� � � �� �� r                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  