pBAV       ��  �� 	  @  ����	�:@   ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  �:    ��������  5F      �����_   � � � �   |5F      �����_   � � � �   @;j$$      �����   � � � �   7j        �����   � � � �   |7         �����   � � � �   @4       �����   � � � �   @@ ((      �����   � � � �   @D ,,      �����   � � � �   @H 00      �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   � z� �F���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              