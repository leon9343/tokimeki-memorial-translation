pBAV       @W ��
   z?  ����.�?   ��������.�?   ��������.�?   ��������.�?   ��������.�?   ��������.�?   ��������.�?   ��������.�?   ��������.�?   ��������.�?   ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    �������� u@5 22      �����_   � � � �  u@2 33      ������   � � � �  J1 //      ������   � � � �  <6 00      ������   � � � �  ,? 11      ������   � � � �  ^R+ )*      ������   � � � �  bR+ ++      ������   � � � �  aR, --      ������   � � � � e,& &&      ������   � � � � eT# $$      ������   � � � �  n@7<<      ������   � � � � @> >>      ������   � � � �  }$? ??      ������   � � � � u@<==      ������   � � � �               ��        � � � �               ��        � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I       ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dx       ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @D       ��ɀ-�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,7        ����-�  � � � � T7        ����-�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @D       ��ɀ-�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dn       ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @=<       ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �   ,��� �F�	:*\��F�@v� N�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        