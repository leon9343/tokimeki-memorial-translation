pBAV        � �� "  x@  ����Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������Ff@   ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������  Ff    ��������@$ $$      ��Ѐ�_   � � � � @& &&      �����_   � � � � 5 55      ��Р�_   � � � � r555      ��Л�_   � � � � n7_ __      �����_   � � � � Z7` ``      �����_   � � � � "0 ++      �����_   � � � � dJ6 66      �����_   � � � � d67 77      �����_   � � � � ^2 ((      �����_   � � � � P"8 88      ����_   � � � � Ph9 99      ����_   � � � � P* **      �����   � � � � K. ..      ��Ѐ�_   � � � � d@# %%      �����_   � � � �               ��        � � � � C        �����_  � � � � hC       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H  L    ����_  � � � � @O M    ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � H        ����_ 	 � � � � |H       ����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,< :@      �����_ 
 � � � � @C AE      �����_  � � � � TH F      �����_  � � � � 7  9      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$  ;    ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  ^F       �����_  � � � �  |^F       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � H        �����_	 	 � � � � |H       �����_	 	 � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �  n@C        �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � P@C       ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   D�4� |�|�P�Tf\�� � ���6 ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                            