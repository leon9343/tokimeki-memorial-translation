pBAV       `�  ��   @  �����@   ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   @< $$      �����   � � � �   @@ ((      �����   � � � �   @D ,,      �����   � � � �   @H 00      �����   � � � �   @L 44      �����   � � � �   @P 88      �����   � � � �   @T <<      �����  	 � � � �   @U @@      �����  
 � � � �   @Q DD      �����   � � � �   @` HH      �����   � � � �   @d LL      �����   � � � �               ��        � � � �               ��        � � � �   �Jd� � � ��.l T��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                