pBAV       0� ��
   o@  ����x ?   ��������d ?   ��������Z ?   ��������Z ?   ��������Z ?   ��������Z ?   ��������Z ?   ��������Z ?   ��������Z ?   ��������Z ?   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������~?& $$      �����_   � � � � ~?% &&      �����_   � � � � ~^7 ))      �����_   � � � � ~O3 --      �����_   � � � � ~(0 //      �����_   � � � � ~/ 22      �����_   � � � � ~61 11      �����_   � � � � ~Z4 33      �����_   � � � � ~?3 44      �����_   � � � � x?4 ::      ��� �_   � � � � ~Z8 88      ��� L   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �  ~?)     ��� �_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?;      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ?Fx     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?T        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ?Pi     ����l�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ?<      ��      � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?DP     ��      � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?C      ��� �_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � d?C      ��� N_	 
 � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �   v���	�lH(��P� �H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                