pBAV       � ��   m@  ����M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������"* **      �����_   � � � � ". ..      �����_   � � � � ", ,,      �����_   � � � � ^7 ))      �����_   � � � � O3 --      �����_   � � � � (0 //      �����_   � � � � / 22      �����_   � � � � 61 11      �����_   � � � � Z4 33      �����_   � � � � @3 44      �����_   � � � � ^5 55      �����_   � � � � @/j$$      ������   � � � � n@3j&&      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � � JTU    ������  � � � � J< T    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O      ����j� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  6H       ������ 	 � � � �  JH       ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @_<S    ��Ȁ��  � � � � @;@ ;      ������  � � � � @w(T    ��Ȁ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @A|     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,T"U    ������  � � � � ,<" T    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ��F��	~*� ~xvF
�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              