pBAV        � ��   @  ����  @   ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������
 @          �����   � � � � 
 @       �����   � � � � 
 @       �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   �#��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        