pBAV       �T �� 0 " l@  ������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    �������� @- $$      ������   � � � � @& &&      ������   � � � �  (* **      ������   � � � �  (, ,,      ������   � � � �  (. ..      ������   � � � � 4 --      ������   � � � � d: ))      ������   � � � � Z7F11      ������   � � � � -7 66      �����_   � � � � <> >>      �����_  	 � � � � F? ??      �����_  
 � � � � P@ @@      �����_   � � � � AD DD      �����_   � � � � U< CC      �����_   � � � � KK KK      ��Ѐ�_   � � � � @U UU      ��Ѐ�_   � � � � 2<  @    ��Ѐ�_  � � � � 2C AE    ��Ѐ�_  � � � � 2H F    ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H H      ��Ѐ�_  � � � � u<
<G      ��Ѐ�_  � � � � k|00;      ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  $      �����_  � � � �   r$     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C  G    ��Ԁ�_  � � � � O H    ��Ԁ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 6<  @      ��Ѐ�_  � � � � JC A      ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n@C      ����_ " � � � � F^C     �����_ " � � � � 2"C     �����_ " � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 7<  @    ��O	  � � � � 7C AE    ��O	  � � � � 7H F    ��O	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � d< @    �����_
  � � � � dCAE    �����_
  � � � � dHF    �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � ZhC
 G    ��Ԁ�_  � � � � ZhO
H    ��Ԁ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 27  9      �����_  � � � � << :@      �����_  � � � � FC AF      �����_  � � � � PH G      �����_   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @ &&      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,H      �����_ ! � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � P@C     ����_ " � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b��� �  �� v 
p \f T F< �r b ~ �J�	�n4 6                                                                                                                                                                                                                                                                                                                                                                                                                                                           