pBAV       @�  ��   @  ����r,@   ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  r,    ��������  @5F      ����P   � � � �   a@4       �����_   � � � �   @8         �����_   � � � �   @< $$      ����@Q   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   �
�$b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      