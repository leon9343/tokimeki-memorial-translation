pBAV       P� �� 	  r@  ����B�@   ��������B�@   ��������B�@   ��������B�@   ��������B�@   ��������B�@   ��������B�@   ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    �������� @)     �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @F:     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � Pi     ������  � � � � rP_     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 7 ,,      ������  � � � � |9d--      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   H�b�
#                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  