pBAV       �� �� -   i@  �����b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������@- $$      ������   � � � � @0 &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ��Ѐ��   � � � � F? ??      ������   � � � � P@ @@      ������   � � � � @% %%      ��Ѐ��   � � � � PA <<      ������   � � � � <> >>      ������   � � � � (I II      ��Ѐ��   � � � � @U UU      ������   � � � � 7<  @    ������ 	 � � � � 7C A    ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C        ������  � � � � |C       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � s
H        �����_  � � � � duH       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � nH        ������  � � � � nl<
       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,[ =      ������  � � � � TC <      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 6<      ����_  � � � � dJ<     �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @+        ��Ѐ�_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @C        �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � I<  @    �����_ 	 � � � � IC A    �����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  YF       �����_  � � � �  rYF       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  YF      �����_  � � � �  rY       �����_  � � � � @0       �����_  � � � � @1       �����_   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 2A<<      ������  � � � � d>>>      ������  � � � � PIII      ��Ѐ��  � � � � d=(==      ������  � � � � ?<??      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,� b��� ��^4*\| �� � � XT��
� < ���b��                                                                                                                                                                                                                                                                                                                                                                                                                                                               