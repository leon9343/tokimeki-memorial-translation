pBAV       ��  ��   @  ����H�@   ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  H�    ��������  @9F      �����   � � � �  6F      �����_   � � � �  r6       �����_   � � � �   |8         �����_   � � � �   8F        �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        