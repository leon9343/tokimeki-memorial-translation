pBAV       �� ��   @  ����  @   ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������  @       �����_   � � � �   @       �����_   � � � �   @(         �����   � � � �   @( $$      �����   � � � �   @< ((      �����   � � � �   @0 ,,      �����   � � � �   @4 00      �����   � � � �   @L 44      �����   � � � �   @F 88      �����  	 � � � �   @P <<      �����  
 � � � �   @L @@      �����   � � � �   @R DD      �����_   � � � �   @Z HH      �����_   � � � �  @\ LL      ��݌�_   � � � �               ��        � � � �               ��        � � � �   �*�� p `�\ � � �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   