pBAV        U  ��   @  ����r�?   ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  @5F      ���� O   � � � �   @3j      �����   � � � �   @=F        �����   � � � �   @>j$$      �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   �\�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      