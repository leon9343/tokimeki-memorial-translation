pBAV       �@ ��   w?  ����d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������d.�@   ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������@Q     �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @O     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � P@Dx     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @8     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Fx9    �����_  � � � � P.x '    �����_  � � � � 2.x(,    �����_  � � � � J.x-8    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @G(     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @.        �����M  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � u3 11      ������  � � � � @0 $$      �����_ 	 � � � � sJ& &&      �����_ 
 � � � � 2 33      ��ʚ-�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @F:       �����M  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<       ����
O	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @I{     �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @5| /      �����_  � � � � f^MT0G      �����_  � � � � M"ehG      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @G( G      �����_  � � � � kkH_      �����_  � � � � Wh�`      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 6Ig     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   X�(����>�\Hvb                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                