pBAV       ��  ��   @  ����  @   ��������  @   ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   @< $$      �����   � � � �   @@ ((      �����   � � � �   @D ,,      �����   � � � �   @H 00      �����   � � � �   @L 44      �����   � � � �   @P 88      �����   � � � �   @T <<      �����  	 � � � �   @X @@      �����  
 � � � �   @\ DD      �����   � � � �   @` HH      �����   � � � �   @d LL      �����   � � � �   @h PP      �����   � � � �   @s TT      �����   � � � �   @4       �����  � � � �   n@3         �����  � � � �   @< $$      �����  � � � �   @?F      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   � �R �� B� � "� � z Rj��� � 8z �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    