pBAV       �� ��   p@  �����b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������d@$ $$      �����_   � � � � d@% &&      �����_   � � � � "* **      �����_   � � � � ". ..      �����_   � � � � ", ,,      �����_   � � � � ^7 ))      �����_   � � � � O3 --      �����_   � � � � (0 //      �����_   � � � � / 22      �����_   � � � � 61 11      �����_   � � � � Z4 33      �����_   � � � � @3 44      �����_   � � � � ^5 55      �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � � @O        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @ID `      ��Ԁ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @)     �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I{     ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Dv       ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ��F��	~H�H�� "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  