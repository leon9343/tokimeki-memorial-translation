pBAV       �z �� ; # s@  ����W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������W�@   ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������  W�    ��������@$ $$      ������   � � � � @# &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))    ������   � � � � Z7F11      ������   � � � � -7 66      ������   � � � � KK KK      ��Ѐ��  	 � � � � @8 88      ��Ѐ��   � � � � KS SS      ������   � � � � nTPTT      �����   � � � � xT
TT      ������   � � � � ^R RR      ��Ѐ��    � � � � n@+  0      ��Ѐ�� 
 � � � � n@7 1D      ��Ѐ��  � � � � dO
EV      ������ 
 � � � � d[
W      ��Д��  � � � � d|OEV      ����� 
 � � � � d|[W      ��Ш��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � d+  -      ��Ѐ��  � � � � d0 .=      ��Ѐ��  � � � � drO>V      ��Ѐ��  � � � � drTW      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � dH        �����  � � � � ,C        �����  � � � � dTO        ������ # � � � � dhH       �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n@<  C      ������  � � � � n@H DK      ������  � � � � @l L      ��Ѐ�� ! � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @$  4      ������  � � � �  d@C 5      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @7  9      ��Ѐ��  � � � � @< :@      ��Ѐ��  � � � � @C A      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n,+  B    ������	  � � � � ndOC    �����	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @C        ������
  � � � � @C        ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � hH E      ������  � � � � $ D      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @+  6    ������  � � � � n@C 7    ����� # � � � � Z^C7    ����� # � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @0  <      ������  � � � � @H =      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � YF@@      ������  � � � � rX @@      ������  � � � � S SS      ������  � � � � n|TTT      ������  � � � � ZF <<      ������ " � � � � ZrF<<      ������ " � � � � d"RRR      ��Ѐ��   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b��� v �F*�.X����^� p � � 4 �	n� ^��f �6                                                                                                                                                                                                                                                                                                                                                                                                                                                         