pBAV       `� ��   i@  ����
M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � -7 66      ������   � � � � @       ��Ѐ��   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �  @$        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � hT R      ������ 	 � � � � @HAQ      ������ 	 � � � � < @      ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @7      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H      ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � "7  ?      ������  � � � � @C @P      ������  � � � � ^O Q      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��Т��	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @<  C      ������
  � � � � @H D      ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �  YF       �����_  � � � �  rYF       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H
       ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� ��� L (\�
"T,l�	n��j @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  