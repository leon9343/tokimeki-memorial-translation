pBAV       �� ��   n?  ����<?   ��������<?   �������� <?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������@5 22      ������   � � � � @3 33      ������   � � � � T1 //      ������   � � � � <6 00      ������   � � � � ,? 11      ������   � � � � %P&&      ����-�  	 � � � � b# $$      ����-�  	 � � � � ^6$P%%      ��ڀ,�  	 � � � � <# ""      ����-�  	 � � � � D! ""      ����-�  	 � � � � @4 44      ������   � � � � Q0 55      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @D     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @+      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��Ɋk�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @A       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @G0       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @R       ��ɀk�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @E     $$��ɀh�	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @P     $$������
 
 � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @"       ������  � � � � @.&&      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @D       �����L  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Dx       ��ۊ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @D       ��ۀ�O  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �Z� Hv����X�	>��6
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            