pBAV       0� ��   |@  ����~�l?   ��������~�l?   ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    ��������  �l    �������� x?&       ��� �_   � � � � 
 ~?2       ��� �_   � � � � 
 v?6         ��� �_   � � � � 
 v?: $$      ��� �_   � � � � 
 v?: ((      ��� �_   � � � � 
 v?= ,,      ��� �_   � � � � 
 z?E 00      ��� �_   � � � � 
 z?H 44      ��� �_   � � � �  d?J 88      ��� �_   � � � �  \?N <<      ��� �_   � � � � 
 p?R @@      ��� �_   � � � �  p?X DD      ��� �_   � � � � 
 p?^ HH      ��� �_   � � � � 
 ~?j LL      ��� �_   � � � �  p?j PP      ��� �_   � � � � 
 d?d TT      ��� �_   � � � �  ~?2       ��� �_  � � � � 
F@3       ��� �_  � � � �  p
6        ��� �_ 	 � � � �  px6<        ��� �_ 	 � � � � X@6 $$      ��� �_ 
 � � � � 
@N((      ��� �_  � � � � 

F((      ��� �_  � � � � 
nF<((      ��� �_  � � � � p?: ,,      ��� �O 
 � � � � p> 00      ���"�M  � � � � pn>00      ��� �M  � � � � l0< 44      ��� �_  � � � � 
?T 88      ��� �_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �ZT�@lv�<���D��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      