pBAV       �� �� D % o@  ����8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������
8@   ��������8@   ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������F7  <    ��Ѐ�_   � � � � FC =    ��Ѐ�_   � � � � d7 <    ��П�_   � � � � dC=    ��П�_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � <7  9      ��ЀJP  � � � � P< :@      ��ЀJP  � � � � dC A      ��ЀJP  � � � � Z27 9      ���JV  � � � � Z<:@      ���JV  � � � � Z
CA      ���JV  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @0      ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$ $$      ��Ѐ�_  � � � �  2& &&      ��Ѐ�_  � � � � 2( ((      �����_  � � � � -* **      �����_ 
 � � � � -, ,,      ��Ѐ�_  � � � � -. ..      ��Ѐ�_  � � � � @3 33      �����_  � � � � (0 00      ��Ѐ�_  � � � � @1 --      ��Ѐ�_  � � � � P2 ))      ��Ѐ�_  � � � � d' ''      �����_ 	 � � � � 2% %%      �����_  � � � � 7? ??      �����_  � � � � 7< @@      �����_  � � � � @0 ##      �����_  � � � �               ��       � � � �  @+      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H      ����IT  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @<        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<  @    ����_  � � � � @C AE    ����_  � � � � @H F    ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � J? CC      �����_  � � � � k"@ DD      �����_  � � � � WTA EE      �����_  � � � � CB FF      �����_  � � � � k?ZCC      ����_  � � � � Wr@ZDD      ����_  � � � � CAZEE      ����_  � � � � /rBZFF      ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$      �����_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �  @H        �����_
 # � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  d@$ $$      �����_ % � � � �        ��Ѐ�_  � � � �        �����_  � � � � ,       �����_  � � � � T       �����_   � � � � P@2 $$      �����_  � � � � @" &&      �����_  � � � � 2* &&      �����_ $ � � � � @       ��Ѐ�_  � � � � h       ��Ѐ�_  � � � � P* **      �����_ " � � � �  dF! ((      �����_ $ � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � YF       �����_ ! � � � � rY        �����_ ! � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  0 <<      �����_  � � � �  1==      �����_  � � � �  "22>>      �����_  � � � �  ,3K??      �����_  � � � �  63 @@      �����_  � � � �  @4AA      �����_  � � � �  J5KBB      �����_  � � � �  T6dCC      �����_  � � � �  ^6DD      �����_  � � � �  h72EE      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @<       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �^� f T �� �	�.
| �� � r b ~ �4 ��� ,�j LNR� *�                                                                                                                                                                                                                                                                                                                                                                                                                                                    