pBAV       �{ ��   s?  ����6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������6L?   ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������  6L    ��������FF 99      ����W   � � � � 8; <<      �����_   � � � � @D DD      ����   � � � �   <F      �����_   � � � �  <F      �����_   � � � � @       �����   � � � �   7       �����   � � � �  7       �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @F     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   <x,6      ������  � � � �  ?<x7<      ������  � � � �  <x=A      ������  � � � � @P Bc      ������  � � � � @"+      ����� 	 � � � �  p dn      ������ 
 � � � � p o      ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <  S    ��      � � � � @dT      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � d< S    �����  � � � � @d
T      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   <        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  <       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<     ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @?m       ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �   �$���� X	~��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     