pBAV       Ф �� 9 , z@  ����8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z;F35      ������   � � � � -7 66      ������   � � � � > >>      ������  	 � � � � <? ??      ������  
 � � � � d@ @@      ������   � � � � (2F12      ������   � � � �               ��        � � � �               ��        � � � � @H AL    �����_  � � � � @O M    ����_  � � � � @0  4    ����_  � � � � @7 5@    ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$  /    ��Ѓ
@  � � � �  @0 0    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � F<      ����_  � � � � n<     ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n,+  +    ��Ѐ�_  � � � � d@0 ,:    ��Ѐ�_  � � � � hO C    ��Ѐ�_  � � � � dT< ;B    ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � JH        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O      ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H K    �����_  � � � � @OL    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � P6H        ����_  � � � � PJ<
       ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T      �����_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � d6$        �����
  � � � � x@$        ����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �  YF<<      �����_  � � � �  |YF<<      �����_  � � � �  5F      �����_  � � � �  T7F      �����_  � � � �  @9F      �����_  � � � �  6:F      �����_   � � � �  
<F      �����_ ! � � � �  P>F!!      �����_ " � � � �  c@F##      �����_ # � � � �  -BF$$      �����_ $ � � � �  ICF&&      �����_ % � � � �  ZEF((      �����_ & � � � �  nGF))      �����_ ' � � � �  PIF++      �����_ ( � � � �               ��       � � � �               ��       � � � � @C      ����,�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,0  9      ������  � � � � @< :G      ������  � � � � TH H      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 5F      �����_ ) � � � � 67F      �����_ * � � � � h9F      �����_ + � � � � |:F      �����_ , � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b��� �  �� � \� ��^*� �|�� ���Vl � � � � � � p � P B ( �                                                                                                                                                                                                                                                                                                                                                                                                                                      