pBAV       � ��
   t@  ����7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������@& $$      �����_   � � � � "* **      �����_   � � � � ". ..      �����_   � � � � ", ,,      �����_   � � � � ^7 ))      �����_   � � � � O3 --      �����_   � � � � (0 //      �����_   � � � � / 22      �����_   � � � � 61 11      �����_   � � � � Z4 33      �����_   � � � � @3 44      �����_   � � � � ^5 55      �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � d@C      ���g�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I       ����*�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C     ��倭� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ���  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @)     ����� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n(I{E    ������  � � � � XI{ D    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C     ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C     ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I        ����*�	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �   v��F��	~��HH� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    