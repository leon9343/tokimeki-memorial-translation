pBAV       �k ��   @  ����8@   ��������
8@   ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  @5F      �����   � � � �   @9F      �����   � � � �   @=F        �����   � � � �   @AF$$      �����   � � � �   @EF((      �����   � � � �   @IF,,      �����   � � � �   @MF00      �����   � � � �   @QF00      �����   � � � �   @QF44      �����   � � � �   @UF88      �����   � � � �   @YF<<      �����  	 � � � �   @]F@@      �����  
 � � � �   @aFDD      �����   � � � �   @eFHH      �����   � � � �   @iFLL      �����   � � � �   @mFPP      �����   � � � �   @5F      �����  � � � �   @<F      �����  � � � �   @=         �����  � � � �   @AF$$      �����  � � � �   @EF((      �����  � � � �   @IF,,      �����  � � � �   @MF00      �����  � � � �   @QF44      �����  � � � �   @UF88      �����  � � � �   @` <<      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   � 2� � 0r.������ ����x� n l NB                                                                                                                                                                                                                                                                                                                                                                                                                                                                                