pBAV        r  ��   @  ����hl?   ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  @0       �����   � � � �   @4       �����   � � � �   @+j        �����   � � � �   @;j$$      �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   �&��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      