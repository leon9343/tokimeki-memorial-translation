pBAV        �  ��   ?  ����.�?   ��������.�?   ��������.�?   ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������@<        ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � mT W      ������  � � � � dT UV      ������  � � � � [T ST      ������  � � � � RT QR      ������  � � � � IT OP      ������  � � � � x@H MN      ������  � � � � x7H KL      ������  � � � � x.H IJ      ������  � � � � x%H GH      ������  � � � � xH DF      ������  � � � � x<  C      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � nT W      ������  � � � � fT UV      ��� ��  � � � � `T ST      ��� ��  � � � � XT QR      ������  � � � � PT OP      ������  � � � � }HH MN      ������  � � � � |@H KL      ������  � � � � {8H IJ      ������  � � � � z0H GH      ������  � � � � y(H EF      ������  � � � � x <  D      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   	"	�	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        