pBAV       � ��   l?  ����@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������@�?   ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    ��������  @�    �������� h@0 22      �����_   � � � � @2 33      ������   � � � � J1 //      ������   � � � � <6 00      ������   � � � � ,? 11      ������   � � � � ]R+ )*      ������   � � � � eR+ ++      ������   � � � � cR, --      ������   � � � � f(& &&      ������   � � � � fX" $$      ������   � � � � J"( ((      ������   � � � �               ������    � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @D       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dx     ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @;.       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T       �����N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @5        ��ڀO  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @D       ��ɀ-�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dy       ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @U s      �����N	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @<       ��7�M
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @I       ��C�N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<
       ��۠JP  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dn     ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I       ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<       ��� j�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   v����F�	:*\x�H�.\�~                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          