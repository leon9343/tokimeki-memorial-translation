pBAV       �� ��   @  ����@   ��������@   ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������      ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   @< $$      �����   � � � �   @< ((      �����   � � � �   @D ,,      �����   � � � �   @H 00      �����   � � � �   @L 44      �����   � � � �   @P 88      �����   � � � �   @T <<      �����   � � � �   @d @@      �����  	 � � � �   @\ DD      �����  
 � � � �   @` HH      �����   � � � �   @d LL      �����   � � � �   @h PP      �����   � � � �   @l TT      �����   � � � �   @8       �����  � � � �   @4       �����  � � � �   @8         �����  � � � �   @D ,,      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �Jdr.l v^ 8JF"�f��N �8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       