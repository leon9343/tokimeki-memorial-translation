pBAV       �K �� '  l@  ����7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������7�@   ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������  7�    ��������@- $$      ������   � � � � @$ &&      ������   � � � � (* **      ������   � � � �  (, ,,      ������   � � � �  (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � -7 66      ������   � � � � Z7 77      ����+�   � � � � @       ������   � � � � P4 44      ��Ѐ+�   � � � � @3j((      ������   � � � � @' ''      ������   � � � �               ��        � � � � @C  E    �����_  � � � � @H F    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ^O 8    ��Ѐ�_ 	 � � � � "C
 7    ��Ѐ�_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$      ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @7      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  H =      ��Ѐ��  � � � �  h$  <      ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @+        ��Ѐ@	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � ,H  C    �����_
  � � � � ZTC     �����_
  � � � � ,T D    �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @<  @    �����_  � � � � @H H    �����_  � � � � @C AG    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @+       ��Ѐ@  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C
       �����_  � � � � rC       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C       �����_  � � � � rC(       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   � b��� f�"x,�
@|\\�r .j �b~ b                                                                                                                                                                                                                                                                                                                                                                                                                                                                         