pBAV        � ��   e@  ����r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������r�@   ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������  r�    ��������@E        �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @O        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dn       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @8        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @7        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ��؀�N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @:        ����O	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @H      �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @4        �����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H =      ���
H 
 � � � � @<  <      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   XX� 2F�Hvb�(�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                