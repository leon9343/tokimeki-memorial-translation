pBAV       �� ��   n@  �����b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������@- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � U' ''      ������   � � � � d2( &&      ��Ѐ��   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � <H  L    ������ 	 � � � � <O M    �����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,7  9      ������  � � � � @< :@      ������  � � � � TC A      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  n@$        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � H :@      ������  � � � � O A      �����_  � � � � C  9      �����_  � � � � hH:@      ������  � � � � hOA      �����_  � � � � hC 9      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � H      �����  � � � � |H     �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C  F    �����  � � � � H G    �����  � � � � |C F    �����  � � � � |HG    �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @P       ����P  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b���� � � f T \�^� �X6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  