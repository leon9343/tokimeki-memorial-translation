pBAV       �
 ��   |@  ����~<?   ��������	~<?   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������
 x?$       ��� �_   � � � � ~
D      ��� �_   � � � � ~nD<      ��� �_   � � � �  z
M        ��� �_   � � � �  ~nM<        ��� �_   � � � � 
Z?D $$      ��       � � � � 
 z?: ((      ��� �_   � � � � 
 z?D ,,      ��� �_   � � � � L?F 00      ��      
 � � � �  ~?P 44      ��       � � � �  f?N 88      ��       � � � �  d?T <<      ��       � � � � 
 ~?\ @@      ��       � � � � 
 ~?h DD      ��      	 � � � � 
 ~?Z HH      ��� �_  	 � � � � 
 ~?X LL      ��� �_   � � � �  ~
F      ��� �_  � � � �  ~xF<      ��� �_  � � � � 
 n(C       ��� �_  � � � � 
 nPB       ��� �_  � � � � 
 ~(=         ��� �_ 	 � � � � 
 ~P>P        ��� �_ 	 � � � � 
 ~??(        ��� �_ 	 � � � � 
 d(J$$      ��� �_  � � � � 
 dPJ
$$      ��� �_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   � �xt�Jzj� ��(4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  