pBAV       �� ��   @  ����y�@   ��������y�@   ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������  y�    ��������?@.C      �����_   � � � � L@4       �����_   � � � � ?@6C        �����_   � � � �  6@:C$$      �����_   � � � � p@@ ((      �����_   � � � � @BC,,      �����_   � � � � |@FC00      �����_   � � � � H@JC44      �����_   � � � � e@NC88      �����_  	 � � � � X@RC<<      �����_  
 � � � �  F@L @@      �����   � � � �  {@\ DD      �����_   � � � �  {@` HH      �����   � � � �   @bCLL      ��� ��   � � � �   @fCPP      ��� ��   � � � �   @jCTT      ��� ��   � � � �  ~@&T      ������  � � � �  }@*T      ������  � � � �  }@.T        ������  � � � �  @2T$$      �����_  � � � �  z@6T((      �����_  � � � �  @:T,,      �����_  � � � �  }@>T00      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ��Z@2R� �������tB�h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      