pBAV       �� ��  	 @  ����	<@   ��������	<@   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������w0  0      ��ݓ�_   � � � � x4 14      ��ݓ�_   � � � � y*7 57      ��ݓ�_   � � � � z5< 8<      ��ݓ�_   � � � � {@@ =@      ��ݓ�_   � � � � |KC AC      ��ݓ�_   � � � � }VH DH      ��ݓ�_   � � � � ~aL IL      ��ݓ�_   � � � � lO M      ��ݓ�_  	 � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � wl0
 0      ��ݓ�_  � � � � xa4
14      ��ݓ�_  � � � � yV7
57      ��ݓ�_  � � � � zK<
8<      ��ݓ�_  � � � � {@@
=@      ��ݓ�_  � � � � |5C
AC      ��ݓ�_  � � � � }*H
DH      ��ݓ�_  � � � � ~L
IL      ��ݓ�_  � � � � O M      ��ݓ�_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ���������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            