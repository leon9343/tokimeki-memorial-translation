pBAV       ��  �� 	 
 q@  ����M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������TC A      ��Ѐ��   � � � � ,<  @      ��Ѐ��   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � 60
     �����  � � � � J<      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � hC        ����_  � � � � @H       ��Ч�_ 	 � � � � O       ��Т�_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   Hbr�� X|�|                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          