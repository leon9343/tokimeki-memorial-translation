pBAV       �� ��   x@  ����n<@   ��������<@   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������d@7  =      ����n�   � � � � d@C >I      ������   � � � � d@O J      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @[        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  d@1 22      ����-�  � � � � @= 33      �����_  � � � � T1 //      �����_  � � � � <6 00      ������  � � � � )? 11      ������  � � � � ^T) )*      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I�      ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @<        ����)� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ����)� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @1       ��ɀ-�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @BF       ����f�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @Uw       ��؀-�	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �  @U       ��؀-�
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �  @C     ��ڀ(�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @;(       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @;       ��      � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @I�       ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � PI�      ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   >�
>�v����4��b.�x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              