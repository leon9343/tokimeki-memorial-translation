pBAV       �� ��   @  ����d@   ��������d@   ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  d    ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   @< $$      �����   � � � �   @< ((      �����   � � � �   @D ,,      �����   � � � �   @H 00      �����   � � � �   @L 44      �����   � � � �   @P 88      �����   � � � �   @T <<      �����   � � � �   @d @@      �����  	 � � � �   @\ DD      �����  
 � � � �   @` HH      �����   � � � �   @d LL      �����   � � � �   @h PP      �����   � � � �   @l TT      �����   � � � �   @0       �����  � � � �   @4       �����  � � � �   @8         �����  � � � �   @< $$      �����  � � � �   @@ ((      �����  � � � �   @D ,,      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �Jdr.l v^ 8JF"�F�z� � N � �8                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   