pBAV       � �� 8  m@  ����M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � AD DD      ������   � � � � U< CC      ������   � � � � KK KK      ��Ѐ��   � � � � @T TT      ������   � � � � @< <<      ������   � � � � @? ??      ������   � � � � @> >>      ������   � � � � @I ==      ������   � � � �  7T @L    ������ 	 � � � �  7[ M    �����_ 
 � � � � d0
 3    ����_ 	 � � � � Z7
4@    ����_ 
 � � � � Z~0 3    ����_ 	 � � � � Z~74@    ����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C  E      �����_  � � � � H F      �����_  � � � � lC E      �����_  � � � � vHF      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � T        �����  � � � � rT       �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 7C        �����_  � � � � dC       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � nH <      �����_  � � � � nH2<      �����_  � � � � nh$  ;      �����_  � � � � nd$2 ;      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � r$  ;    ����_  � � � � 0 ;    ����_  � � � � O <      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 2C  L      �����_	  � � � � NOM      �����_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � 6H        ����_
  � � � � d@C        ����_
  � � � � dJH       ����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � 6H =T    �����_  � � � � 6T U    �����_  � � � � FJ0
 6    ����_  � � � � FJ<
7<    ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n<<        �����_  � � � � d@<(       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C      ����_  � � � � rC     ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <        �����_  � � � � r<
       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � n@C        �����_  � � � � n@<
       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �� ���� v < � � �\.J�
�� � p �Fr ~ �	4��*�                                                                                                                                                                                                                                                                                                                                                                                                                                                                