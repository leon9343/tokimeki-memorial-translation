pBAV       �) ��   i@  ����B�@   ��������B�@   ��������B�@   ��������B�@   ��������B�@   ��������B�@   ��������B�@   ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������  B�    ��������@& $$      ������   � � � � @% &&      ������   � � � � "* **      ������   � � � � ". ..      ������   � � � � ", ,,      ������   � � � � ^7 ))      ������   � � � � O3 --      ������   � � � � (0 //      ������   � � � � / 22      ������   � � � � 61 11      ������   � � � � Z4 33      ������   � � � � @3 44      ������   � � � � ^5 55      ������   � � � � EA 66      �����_    � � � � <7 77      �����_    � � � �               ��        � � � �  @+      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      ���i�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @_<S    ��Ȁ�� 	 � � � � @;@ ;      ������ 
 � � � � @w(T    ��Ȁ�� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @O
N      ����*�  � � � � @Dx M      ����*�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dv       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   v���F��	~~x2��b ��4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            