pBAV        � �� -   j@  ������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������@   ����������   ����������@   ����������@   ����������@   ��������d��@   ����������@   ����������@   ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    ��������  ��    �������� &  +      ������   � � � �  Z2 ,9      ������   � � � �  ?J CO      ������   � � � �  Z?V P      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �  @< G    �����  � � � �  @[ H    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$ $$      �����  � � � � @& &&      �����  � � � � 
. ))      �����  � � � � @, --      ������  � � � � u* 00      ������  � � � � @% %%      ������  � � � �  d+ ++      ������  � � � � @F HH      �����  � � � � @J JJ      �����  � � � �  @0 ""      ������  � � � � ,<##      ������  � � � � T7m!!      �����  � � � �  
T TT      �����  � � � �  uV VV      �����  � � � �  2X XX      �����  � � � �  TY YY      �����  � � � � ?<  A    �����X  � � � � FbB    ��ˎ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C  S      ����@� 
 � � � � @` T      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � dO <      ����_ 	 � � � � +  ;      ����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  H        ����^�  � � � � ?H       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @< 0     ������  � � � �  <
0     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @7      �����	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @<        �����_
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �  @<        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  F@
 (      ����   � � � �  F9 )P      ����   � � � �  FP Qx      ����   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  nnF=Z      �����_  � � � �  nzFQ      �����_  � � � � @/v <      �����_   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ��ۘ�_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � dx<       ����O_  � � � � d<       ����O  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   h�6�p�X4� D *P<$"���|4 � l� � f"&                                                                                                                                                                                                                                                                                                                                                                                                                                                              