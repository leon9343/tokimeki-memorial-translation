pBAV       �1 ��   @  �����b@   ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������
 @F      �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   �D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            