pBAV       �e ��   g@  ����  @   ��������  @   ��������  @   ��������  @   ��������  @   ��������  @   ��������  @   ��������  @   ��������  @   ��������n  @   ��������  @   ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        �������� d@O  F      ������   � � � �  d@T G      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @7  =      �����  � � � � @C>I      ������  � � � � @OJ      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @7        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<       ����D�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  J[  O      ����� 	 � � � �  6[ P      ����� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � T <      ����� 
 � � � �  0 ;      ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @H        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  J[  O      ����� 	 � � � �  6[ P      ����� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � d@7  =      ����N_	  � � � � d@C >I      �����_	  � � � � d@O J      �����_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @[        ������
 	 � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �   |�.Tp�� >
�
>�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    