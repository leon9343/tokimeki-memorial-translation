pBAV       `�  �� 
  @  ����
8@   ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  @0       �����   � � � �   @4       �����   � � � �   @8         �����   � � � �   @< $$      �����   � � � �   @@ ((      �����   � � � �   @9 ,,      �����   � � � �   @A 00      �����   � � � �   @I 44      �����   � � � �   @Q 88      �����   � � � �   @Y <<      �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   F<T�� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  