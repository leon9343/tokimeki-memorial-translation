pBAV       P�  ��   ?  ����Y�?   ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  Y�    ��������  |@/C      ������   � � � �   |@(       ��ʀ �   � � � �   @=F        ������   � � � �   F: $$      ������   � � � �   :@
((      ������   � � � �   Y@7F,,      �����   � � � �   Z0; ##      ������   � � � �   PFA<((      ������   � � � �               ��        � � � �               �� � �    � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   ��`�N`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   