pBAV       0� ��   w?  ����<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    �������� c@/22      ������   � � � � o@2 33      ������   � � � � iT. //      ������   � � � � k<3&00      ������   � � � � m,< 11      ������   � � � � ^^) ))      ������   � � � � p^+ ++      ������   � � � �  a^- --      ������   � � � � d& &&      ������   � � � � db" $$      ������   � � � � W74 44      ������   � � � � [75 55      ������   � � � � S1 66      �����_   � � � � n^* **      ����,�   � � � �              ������    � � � �               ��        � � � � @D       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @P A      ��ˀ��  � � � � @UB~      ����(� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        �����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Q        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � u@Q        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        �����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        �����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @P C      ������  � � � � @UD~      ������ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @Dy       ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @P       ��� (�
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @5        ��ڔ�O  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   v�����	�6�\.�
XF�H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            