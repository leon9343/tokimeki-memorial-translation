pBAV       Pr ��   @  ����+�@   ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  +�    ��������  @*F      �����   � � � �   @4       �����   � � � �   >F        �����   � � � �   r>F        �����   � � � �   @<F$$      �����   � � � �   HF((      �����   � � � �   rHF((      �����   � � � �   @8 ,,      �����   � � � �   @HF00      �����  	 � � � �   @HF44      �����  
 � � � �   @P 88      �����   � � � �   @T <<      �����   � � � �   @]F@@      �����   � � � �   @aFDD      �����   � � � �   Z@T HH      �����   � � � �               ��        � � � �   �X��r��N�� $����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                