pBAV       @� �� 3  m@  ����o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������o�@   ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������  o�    ��������@- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ��Ѐ��   � � � � 7 66      ��Ѐ��   � � � � Z' ''      ��Ѐ��   � � � � 2K KK      ������   � � � � F< <<      ������   � � � � (> >?      ������   � � � � I II      ��Ѐ��   � � � � @4j((      ������   � � � � 7C AG    �����  � � � � 7<  @    �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � +
     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  6$  ;    ������ 	 � � � � J[ <      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � TC  R    ����� 
 � � � � d[S    ����� 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<  G      ������  � � � � @T
H      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,<  G    ��݀��  � � � � ZJT H    �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C  H    ������  � � � � d[
I      ������  � � � � d|[I      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 6C      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 
<  H      ������	  � � � � vA  H      ������	  � � � � dTI      ������	  � � � � d|YI      ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � x
C        ������
  � � � � Z@H        �����
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � C        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @$  ;    ������  � � � � @> >>      ������  � � � � d?(??      ������  � � � � P|@P@@      ������  � � � � 6A <<      ������  � � � � (I II      ��Ѐ��  � � � � ddJJJ      ��Ч��  � � � � hB ==      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � JH      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ZH        �����  � � � � H       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <        ������  � � � � |<       �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b���b \� � �Xfp B�L  v ��b r �b�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                