pBAV       �+ ��   h@  �����>@   ���������>@   ���������>@   ���������>@   ���������>@   ���������>@   ���������>@   ���������>@   ���������>@   ���������>@   ���������>@   ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    ��������  �>    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � P' ''      ������   � � � � d(D DD      ������   � � � � (K KK      ������   � � � � 7 66      ������   � � � � ZA AA      ������   � � � � d(< CC      ������   � � � � dPDDD      ������   � � � � dP<CC      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � � @<  B      ������  � � � � @C CE      �����_  � � � � @H F      �����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @$        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � "H  L    ������  � � � � "O M    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ^H L    ������	  � � � � ^OM    ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @P       ����P
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �   ,�� b�r b ~ � � \� v  ���|6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      