pBAV       �l  ��   @  ����hl?   ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  hl    ��������  5      �����_   � � � �   r5      �����_   � � � �   @3j      �����_   � � � �   @+j        �����   � � � �   @AF$$      �����   � � � �   @?j((      �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   ��d��n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  