pBAV       �n ��   ~?  ����<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������<?   ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������  <    ��������a74 44      ������   � � � � \73 33      ������   � � � � W72 22      ������   � � � � R71 11      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � @P       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��ɀk�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @A ?      �����N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @F8       ��ր�N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @F8       ��ր�N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H
       ��ɀk�	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @H        ��ɀk�
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @E	       ��ɔHV  � � � �               ��ɨHV   � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @E        ��ɔHV  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @E       ��ɔHV  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   .�6\HvbX                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              