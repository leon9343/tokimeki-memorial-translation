pBAV         �� "  p@  ����M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������M�@   ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    ��������  M�    �������� Gj<<      �����_   � � � � ,Gj>>      �����_   � � � � |G <<      �����_   � � � � dhH??      �����_   � � � � dHj??      �����_   � � � � @$ $$      �����_   � � � � ,& &&      �����_   � � � � ,) ))      �����_   � � � � ,( ((      �����_   � � � � * **      �����_   � � � � . ..      �����_   � � � � J0 00      �����_   � � � � @0j##      �����_   � � � � 9j""      �����_   � � � � |9 ""      �����_   � � � �               ��        � � � � @7        ����
@  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ����@  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <        �����_  � � � � Z|<(       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @J        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � d6C        �����_  � � � � nJ7        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C     �����_  � � � � d|C(     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$        ��Ѐ@ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @+        ��Ѐ@  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,C        ��Ѐ�_	  � � � � TC        ��Ѐ�_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @H      �����_
 
 � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @C      ��Ѐ@  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <       �����_  � � � � d|<       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @J        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @J        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   .Z�� � � � � �XZ� ��	$��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                