pBAV       �� �� "  j@  �����@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ���������@   ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������  �    ��������* **      ������   � � � � . ..      ������   � � � � ^2 ))      ������   � � � � O- --      ������   � � � � <* //      ������   � � � � ( 22      ������   � � � � 0 11      ��Ѐ��   � � � � J2 33      ��Ѐ��   � � � � ^4 44      ��Ѐ��   � � � � T5 55      ������   � � � � s@" &&      ������   � � � � n@& $$      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �  ;=H    ������  � � � �  ;ZFI`    ������  � � � �  ;     ��b���  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @TUf    ������  � � � � @< T    ������  � � � � @lg    �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @_<S    ��Ȁ�� 	 � � � � u@;  ;      ������ 
 � � � � @w(T    ��Ȁ�� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 6<  `    ������  � � � � Jl a    �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C T    ������  � � � � @s`    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @=x T      ��G�c�  � � � � @mxU      ��G�i�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @<     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @F0       ��ʀ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � F0       ��ʀ��	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � F0       ��ʀ��
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @C        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @0        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ���	~@b*~xH��� ,4 ��b                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    