pBAV       � ��    m@  ����Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������Z@   ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������  Z    ��������@- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � d-& &&      ������   � � � � @% %%      ������   � � � � 7 ##      ������   � � � � ^6 ""      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �  @$      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      ������  � � � � nC     �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � C      	�����  � � � � PhC
     	������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � "7  2      ��Ѐ��  � � � � @7 2<      ��Ѐ��  � � � � ^7 =      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  YF<<      �����_  � � � �  drYF<<      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @C        ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ,O        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � dTO
       ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b��� �  �� v �B@f�F���                                                                                                                                                                                                                                                                                                                                                                                                                                                                               