pBAV       0�  ��   n@  ����.�@   ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    �������� |@0       ������   � � � � |@(       ������   � � � � `@8         ������   � � � � |@< $$      ������   � � � � p@>C((      ������   � � � � @D ,,      ������   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   �
���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  