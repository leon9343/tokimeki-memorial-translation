pBAV       ��  ��   @  ����8>@   ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  8>    ��������  @0       �����   � � � �   @;F      �����   � � � �   @=F        �����   � � � �   @Bm$$      �����   � � � �   @?F((      �����   � � � �   @D ,,      �����   � � � �   @H 00      �����   � � � �   @VF44      �����   � � � �   @TF88      �����   � � � �   @VF<<      �����   � � � �   @XF@@      �����   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   ,���� ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              