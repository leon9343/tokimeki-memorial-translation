pBAV       P� ��
   ?  ����  ?   ��������  ?   ��������  ?   ��������  ?   ��������  ?   ��������  ?   ��������  ?   ��������  ?   ��������  ?   ��������  ?   ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        �������� c@5 22      ������   � � � � u@2 33      ������   � � � � J2 //      ������   � � � � <; 00      ������   � � � � ,? 11      ������   � � � � `T) ))      ������   � � � � dT+ ++      ������   � � � � _T- --      ������   � � � � g(& &&      ������   � � � � gX" $$      ������   � � � � T* **      ����,�   � � � � _T. ..      ������   � � � �               ������    � � � �               ������    � � � �               ������    � � � �               ��        � � � � @P       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H       ��ƀ)�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��ɀk�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @5       �����N  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T       �����Q  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @P       ��� (�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H       ��ɀ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��x �^	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �   v������	.�
6\HvF�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              