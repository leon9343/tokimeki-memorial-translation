pBAV       `�  ��   z@  ����.�@   ��������.�@   ��������.�@   ��������.�@   ��������.�@   ��������.�@   ��������.�@   ��������.�@   ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������  .�    ��������
7  9      �����_   � � � � < :@      �����_   � � � � C A      �����_   � � � �  d7 9      ��Ш�_   � � � �  n<:@      ��Ш�_   � � � �  xCA      ��Ш�_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �  @<  @      ��݀�_  � � � �  @C A      ��݀�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @0        ��Ш�_  � � � �  d<
       ����_  � � � �  dr0       ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  <7  9      ��Ѐ�_  � � � �  @< :@      ��Ѐ�_  � � � �  FC A      ��Ѐ�_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @* **      ������ 
 � � � �  @. ..      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  <
 @      �����_  � � � �  C
A      �����_  � � � �  r< @      ����_  � � � �  rCA      ��ݭ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  <7 9      ��Ѐ�_  � � � �  @<:@      ��Ѐ�_  � � � �  FCA      ��Ѐ�_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  C        ����_  � � � �  |C       ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   �rb� � ��VF�	X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      