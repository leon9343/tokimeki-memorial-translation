pBAV       �� ��   t@  ����x ?   ��������V ?   ��������d ?   ��������d ?   ��������d ?   ��������d ?   ��������d ?   ��������d ?   ��������d ?   ��������d ?   ��������d ?   ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������       ��������d?& $$      �����_   � � � � d?% &&      �����_   � � � � d"* **      �����_   � � � � d". ..      �����_   � � � � d^7 ))      �����_   � � � � dO3 --      �����_   � � � � d(0 //      �����_   � � � � d/ 22      �����_   � � � � d61 11      �����_   � � � � dZ4 33      �����_   � � � � d?3 44      �����_   � � � � d^5 55      �����_    � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � d?O      ����j�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?I       ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  ?)     ����� 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?I{       ������ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?Dx       ����+�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � x?T        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~?;        ��� �_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � ~F;       ��� �_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � t?<        ��� �_	  � � � � t?<
       ��� �_	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � x?T        ��    
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �   v�����	� HH��	ZP�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 