pBAV       P� ��    e@  �����b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ���������b@   ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    ��������  �b    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � � (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � -7 66      ������   � � � � KK KK      ��Ѐ��  	 � � � � ,O OO      ����,�  
 � � � � ,N NN      ������   � � � � J' ''      ������   � � � � @4 44      ������   � � � � #( 22      ������   � � � � H        ������  � � � � drH       ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � 7C      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <H      �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  YF       �����_  � � � �  |YF       �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @%( <    ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � JH      ������	  � � � � 6H
     �����	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @C      ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � @7      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @C        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b��� v �.��p � �F��@@�T�
�                                                                                                                                                                                                                                                                                                                                                                                                                                                                         