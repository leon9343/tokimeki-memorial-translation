pBAV       p� ��  
 r@  ����;@@   ��������;@@   ��������;@@   ��������;@@   ��������;@@   ��������;@@   ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������  ;@    ��������+73:    �����_   � � � � +>;A    �����_   � � � � +CBF    �����_   � � � � +JGL    �����_   � � � � +OMS    �����_   � � � � +\T    �����N   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � � S7 3:    �����_  � � � � S> ;A    �����_  � � � � SC BF    �����_  � � � � SJ GL    �����_  � � � � SO MS    �����_  � � � � S\	T    �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @9     ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  <  <    �����  � � � � T=    �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @<        �����_ 	 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @<        �����_ 
 � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   @���4�� �P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          