pBAV        �  ��   P@  ����w^@   ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  w^    ��������  0       �����_   � � � �   |0       �����_   � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �               ��        � � � �   ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          