pBAV        � �� '  p@  ����8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������8@   ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    ��������  8    �������� @- $$      ������   � � � � @& &&      ������   � � � � (* **      ������   � � � � (, ,,      ������   � � � �  (. ..      ������   � � � � (0 00      ������   � � � � @4 --      ������   � � � � P: ))      ������   � � � � Z7F11      ������   � � � � -7 66      ������   � � � � <> >>      ������  	 � � � � F? ??      ������  
 � � � � P@ @@      ������   � � � � AD DD      ������   � � � � U< CC      ������   � � � � KK KK      ��Ѐ��   � � � � @C      ��٣*�  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        �����  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � <7  <    ��Ѐ��  � � � � FC =    ��Ѐ�_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � x
T I      ������  � � � � Z<1H      ��Ѐ��  � � � � F|$
 0      ��Ѐ��  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @O        ����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @H  K      ������  � � � � @O L      ������  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  @$      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @<        �����	  � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � �               ��    	   � � � � @H        ������
  � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � �               ��    
   � � � � ;<  D      ������  � � � � EH E      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @T        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � @$        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � � x<<        �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �  YF<<      �����_  � � � �  rYF<<      �����_  � � � �  [F>>      �����_  � � � �  r[F>>      �����_  � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �               ��       � � � �   ,�� b��� �  �� v � � \� �^*�|��	nlll��                                                                                                                                                                                                                                                                                                                                                                                                                                                                